//`timescale 1 ns/100 ps


module tb_6bit;
 // signal declaration
   reg  [5:0]a,b;
   reg [2:0] fxn;
  
   wire [5:0] OUT;
   wire C,V;
   // instantiate the circuit under test
   main uut
      (.a(a),.b(b), .fxn(fxn),.OUT(OUT),.Cled(C),.Vled(V));

   //  test vector generator
   initial
   begin
   $monitor ("INPUT = %d",a);
   $monitor ("FXN = %d",fxn);
   $monitor ("OUTPUT =  %d",OUT);
   $monitor ("CARRY =%d",C);
   $monitor ("OVERFLOW = %d",V);




    // test vector 1
//      fxn = 3'b000;
//      a = 6'b001100; //First 6 digits of Board number..
//      b =  6'b000001;
//      # 100;
//       a = 6'b000000;
//      b = 6'b000000;
//      # 100;
//      a = 6'b000001; //
//      b = 6'b000001;
//      # 100;
//      a = 6'b100000; //
//      b = 6'b100000;
//      # 100;
//      a = 6'b101010; //
//      b = 6'b101010;
//      # 100;
//      a = 6'b101111; //
//      b = 6'b101010;
//      # 100;
//      a = 6'b101111; //for a<b
//      b = 6'b111111;
//      # 100;
//      a = 6'b101000; //
//      b = 6'b101010;
//      # 100;
    //////////////////////////////
//      // test vector 2//Basic input testing
//      fxn = 3'b001;
//       a = 6'b001100; //First 6 digits of Board number..
//      b =  6'b000001;
//      # 100;
//       a = 6'b000000;
//      b = 6'b000000;
//      # 100;
//      a = 6'b000001; //
//      b = 6'b000001;
//      # 100;
//      a = 6'b100000; //
//      b = 6'b100000;
//      # 100;
//      a = 6'b101010; //
//      b = 6'b101010;
//      # 100;
//      a = 6'b101111; //
//      b = 6'b101010;
//      # 100;
//      a = 6'b101111; //for a<b
//      b = 6'b111111;
//      # 100;
//      a = 6'b101000; //
//      b = 6'b101010;
//      # 100;
//      a = 6'b000000;
//      b =  6'b111111;
//      # 100;
//       ////////////////////////////// -A
         // test vector 2
//      fxn = 3'b010;
//       a = 6'b001100; //First 6 digits of Board number..
//      b =  6'b000001;
//      # 100;
//       a = 6'b000000;
//      b = 6'b000000;
//      # 100;
//      a = 6'b000001; //
//      b = 6'b000001;
//      # 100;
//      a = 6'b100000; //
//      b = 6'b100000;
//      # 100;
//      a = 6'b101010; //
//      b = 6'b101010;
//      # 100;
//      a = 6'b101111; //
//      b = 6'b101010;
//      # 100;
//      a = 6'b101111; //for a<b
//      b = 6'b111111;
//      # 100;
//      a = 6'b101000; //
//      b = 6'b101010;
//      # 100;
//      a = 6'b101010;
//      b =  6'b111111;
//      # 100;
      
//    //////////////////////////////////////-B
//      fxn = 3'b011;
//       a = 6'b001100; //First 6 digits of Board number..
//      b =  6'b000001;
//      # 100;
//       a = 6'b000000;
//      b = 6'b000000;
//      # 100;
//      a = 6'b000001; //
//      b = 6'b000001;
//      # 100;
//      a = 6'b100000; //
//      b = 6'b100000;
//      # 100;
//      a = 6'b101010; //
//      b = 6'b101010;
//      # 100;
//      a = 6'b101111; //
//      b = 6'b101010;
//      # 100;
//      a = 6'b101111; //for a<b
//      b = 6'b111111;
//      # 100;
//      a = 6'b101000; //
//      b = 6'b101010;
//      # 100;
//      a = 6'b101010;
//      b =  6'b101010;
//      # 100;
      
//      /////////////////////////////////// A<B
//         // test vector 2
      fxn = 3'b100;
       a = 6'b001100; //First 6 digits of Board number..
      b =  6'b000001;
      # 100;
       a = 6'b000000;
      b = 6'b000000;
      # 100;
      a = 6'b000001; //
      b = 6'b000001;
      # 100;
      a = 6'b100000; //
      b = 6'b100000;
      # 100;
      a = 6'b101010; //
      b = 6'b101010;
      # 100;
      a = 6'b101111; //
      b = 6'b101010;
      # 100;
      a = 6'b101111; //for a<b
      b = 6'b111111;
      # 100;
      a = 6'b101000; //
      b = 6'b101010;
      # 100;
      a = 6'b101010;
      b =  6'b111111;
      # 100;
      
//      ///////////////////////////////////XNOR
     
//      fxn = 3'b101;
//       a = 6'b001100; //First 6 digits of Board number..
//      b =  6'b000001;
//      # 100;
//       a = 6'b000000;
//      b = 6'b000000;
//      # 100;
//      a = 6'b000001; //
//      b = 6'b000001;
//      # 100;
//      a = 6'b100000; //
//      b = 6'b100000;
//      # 100;
//      a = 6'b101010; //
//      b = 6'b101010;
//      # 100;
//      a = 6'b101111; //
//      b = 6'b101010;
//      # 100;
//      a = 6'b101111; //for a<b
//      b = 6'b111111;
//      # 100;
//      a = 6'b101000; //
//      b = 6'b101010;
//      # 100;
//      a = 6'b101010;
//      b =  6'b111111;
//      # 100;
//      //////////////////////////////////A+B
//      fxn = 3'b110;
//       a = 6'b001100; //First 6 digits of Board number..
//      b =  6'b000001;
//      # 100;
//       a = 6'b000000;
//      b = 6'b000000;
//      # 100;
//      a = 6'b000001; //
//      b = 6'b000001;
//      # 100;
//      a = 6'b100000; //
//      b = 6'b100000;
//      # 100;
//      a = 6'b101010; //
//      b = 6'b101010;
//      # 100;
//      a = 6'b101111; //
//      b = 6'b101010;
//      # 100;
//      a = 6'b101111; //for a<b
//      b = 6'b111111;
//      # 100;
//      a = 6'b101000; //
//      b = 6'b101010;
//      # 100;
//      a = 6'b101010;
//      b =  6'b111111;
//      # 100;
      
//      ///////////////////////////////A-B
      
//        fxn = 3'b111;
//         a = 6'b001100; //First 6 digits of Board number..
//      b =  6'b000001;
//      # 100;
//       a = 6'b000000;
//      b = 6'b000000;
//      # 100;
//      a = 6'b000001; //
//      b = 6'b000001;
//      # 100;
//      a = 6'b100000; //
//      b = 6'b100000;
//      # 100;
//      a = 6'b101010; //
//      b = 6'b101010;
//      # 100;
//      a = 6'b101111; //
//      b = 6'b101010;
//      # 100;
//      a = 6'b101111; //for a<b
//      b = 6'b111111;
//      # 100;
//      a = 6'b101000; //
//      b = 6'b101010;
//      # 100;
//      a = 6'b101010;
//      b =  6'b111111;
//      # 100;
//      fxn = 3'b111;
//      a = 6'b000000;
//      b =  6'b000000;
//      # 100;
      
//      fxn = 3'b111;
//      a = 6'b111000;
//      b =  6'b000111;
//      # 100;
      
//       fxn = 3'b110;
//      a = 6'b111110;
//      b =  6'b110111;
//      # 100;
//      fxn = 3'b110;
//      a = 6'b101010;
//      b =  6'b111111;
//      # 100;
//      fxn = 3'b110;
//      a = 6'b000000;
//      b =  6'b000000;
//      # 100;
      
//      fxn = 3'b110;
//      a = 6'b111000;
//      b =  6'b000111;
//      # 100;
      
//       fxn = 3'b110;
//      a = 6'b111110;
//      b =  6'b110111;
//      # 100;
//        stop simulation
      $stop;
   end
 endmodule
